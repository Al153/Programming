----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:09:43 04/05/2006 
-- Design Name: 
-- Module Name:    sram_interface - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity sram_sm is
    Port ( sm_clk_in : in std_logic;
			  fpga_clk_in : in std_logic;
           rst_in : in std_logic;	 
			  a : out  STD_LOGIC_VECTOR (16 downto 0);
           din : in  STD_LOGIC_VECTOR (7 downto 0);
           dout : out  STD_LOGIC_VECTOR (7 downto 0);
			  dir : out std_logic;
           oe_n : out  STD_LOGIC;
           we_n : out  STD_LOGIC;
			  errors : out  STD_LOGIC_VECTOR (16 downto 0);
			  test_failed : out std_logic);
end sram_sm;

architecture rtl of sram_sm is

   type state_type is (st1_w0_idle, st2_w1_addr, st3_w2_data, st4_w3_hold,
	                    st5_w4_d_en, st6_w5_d_a, st7_r0_idle, st8_r1_addr,
							  st9_r2_oe, st10_r3_hold, st11_r4_data, st12_r5_comp); 
   signal state, next_state : state_type; 

   signal oe_n_int : STD_LOGIC;
   signal we_n_int : STD_LOGIC;
   signal dir_int,dir_copy : STD_LOGIC;
   signal errors_int : STD_LOGIC_VECTOR (16 downto 0);
	signal test_failed_int : STD_LOGIC;
	
   signal count : STD_LOGIC_VECTOR (16 downto 0);
   signal result : STD_LOGIC_VECTOR (7 downto 0);
   signal value : STD_LOGIC_VECTOR (7 downto 0);
   signal reset_count,reset_count_int : std_logic;
   signal increment,store_value,comp_value : std_logic;
   signal increment_int,store_value_int,comp_value_int : std_logic;
	
	signal rst_in_d, rst_in_d2 : std_logic;
	signal start : std_logic; 
	signal start_p : std_logic;

begin

   -- The Edge Detect process detects the falling edge of reset
	-- and creates the state machine state strobe as follows:
	--            ________
	--     rst_in         |__________
	--            __________
	--   rst_in_d           |________
	--            ____________
	--  rst_in_d2             |______
   --                       _
   --    start_p __________| |______	
	--
	edge_detect : process(fpga_clk_in)
	begin
      if (fpga_clk_in'event and fpga_clk_in = '1') then
         rst_in_d <= rst_in; -- rst_in delayed one clock
			rst_in_d2 <= rst_in_d; -- rst_in delayed two clocks
			-- start strobe asserts high one clock on reset deassert
			start_p <= rst_in_d2 AND NOT(rst_in_d); -- reset deassert
			start <= start_p; --add another clock of seperation after reset
		end if;
	end process;	

	-- SRAM test - writes sram with a counting pattern equivalent
	-- to the data values address in memory, reads back the data
	-- written and compares it to the expect value (its address).
	-- The test starts once on reset deassert as generated by the 
	-- Edge Detect process.

   -- The Sram_test_sync Process is the synchronous part of the
	-- Moore state machine 
   sram_test_sync: process (sm_clk_in)
   begin
      if (sm_clk_in'event and sm_clk_in = '1') then
         if (rst_in = '1') then
            state <= st1_w0_idle;
            oe_n 	<= '1'; -- active low
            we_n 	<= '1'; -- active low
				dir 	<= '1'; -- 1 = read, 0 = write (data out enabled)
				dir_copy <= '1'; -- copy of dir for internal use
				store_value <= '0'; -- store data in & expected value
				increment <= '0'; -- increment address counter
				comp_value <= '0'; -- compare data in & expected value
				reset_count <= '1'; -- reset address counter
        else
            state <= next_state;
            oe_n 	<= oe_n_int;
            we_n 	<= we_n_int;
				dir 	<= dir_int;
				dir_copy <= dir_int;
				store_value <= store_value_int;
				increment <= increment_int;
				comp_value <= comp_value_int;
				reset_count <= reset_count_int;
         end if;        
      end if;
   end process;
 
   -- The Sram_test_output_decode Process is the combinatorial output
   -- decode part of the Moore state machine.  
   -- In a MOORE State Machine the outputs are based on the state only
   sram_test_output_decode: process (state)
   begin      
		case (state) is
         when st1_w0_idle =>
            oe_n_int 	<= '1';
            we_n_int 	<= '1';
				dir_int 	<= '1'; -- read (output disabled)
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '1'; --reset address counter
         when st2_w1_addr =>
			-------------------	
			-- Write State 1 --
			-------------------
            oe_n_int 	<= '1';
				------------------------------------------------
            we_n_int 	<=      --** Add write strobe output
				                    --** value for W1 state         
				------------------------------------------------
				dir_int 	<= '0';
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '0';
         when st3_w2_data =>
			-------------------	
			-- Write State 2 --
			-------------------
            oe_n_int 	<= '1';
				------------------------------------------------
            we_n_int 	<=      --** Add write strobe output
				                    --** value for W2 state         
				------------------------------------------------
				dir_int 	<= '0'; -- write (data out enabled)
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '0';
         when st4_w3_hold =>
			-------------------	
			-- Write State 3 --
			-------------------
            oe_n_int 	<= '1';
				------------------------------------------------
            we_n_int 	<=      --** Add write strobe output
				                    --** value for W3 state         
				------------------------------------------------
				dir_int 	<= '0'; -- write (data out enabled)
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '0';
         when st5_w4_d_en =>
			-------------------	
			-- Write State 4 --
			-------------------
            oe_n_int 	<= '1';
				------------------------------------------------
            we_n_int 	<=      --** Add write strobe output
				                    --** value for W4 state         
				------------------------------------------------
				dir_int 	<= '0'; -- write (data out enabled)
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '0';
         when st6_w5_d_a =>
			-------------------	
			-- Write State 5 --
			-------------------
            oe_n_int 	<= '1';
				------------------------------------------------
            we_n_int 	<=      --** Add write strobe output
				                    --** value for W5 state         
				------------------------------------------------
				dir_int 	<= '0'; -- write (data out enabled)
				store_value_int <= '0';
				increment_int <= '1'; -- increment address counter
				comp_value_int <= '0';
				reset_count_int <= '0';
         when st7_r0_idle =>
            oe_n_int 	<= '1';
            we_n_int 	<= '1';
				dir_int 	<= '1'; -- read (output disabled)
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '1'; --reset address counter
         when st8_r1_addr =>
			------------------	
			-- Read State 1 --
			------------------
				------------------------------------------------
            oe_n_int 	<=      --** Add write strobe output
				                    --** value for R1 state         
				------------------------------------------------
            we_n_int 	<= '1';
				dir_int 	<= '1'; -- read (output disabled)
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '0';
         when st9_r2_oe =>
			------------------	
			-- Read State 2 --
			------------------
				------------------------------------------------
            oe_n_int 	<=      --** Add write strobe output
				                    --** value for R2 state         
				------------------------------------------------
            we_n_int 	<= '1';
				dir_int 	<= '1'; -- read (output disabled)
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '0';
         when st10_r3_hold =>
			------------------	
			-- Read State 3 --
			------------------
				------------------------------------------------
            oe_n_int 	<=      --** Add write strobe output
				                    --** value for R3 state         
				------------------------------------------------
            we_n_int 	<= '1';
				dir_int 	<= '1'; -- read (output disabled)
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '0';
         when st11_r4_data =>
			------------------	
			-- Read State 4 --
			------------------
				------------------------------------------------
            oe_n_int 	<=      --** Add write strobe output
				                    --** value for R4 state         
				------------------------------------------------
            we_n_int 	<= '1';
				dir_int 	<= '1'; -- read (output disabled)
				store_value_int <= '1'; -- store read value
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '0';
         when st12_r5_comp =>
			------------------	
			-- Read State 5 --
			------------------
				------------------------------------------------
            oe_n_int 	<=      --** Add write strobe output
				                    --** value for R5 state         
				------------------------------------------------
            we_n_int 	<= '1';
				dir_int 	<= '1'; -- read (output disabled)
				store_value_int <= '0';
				increment_int <= '1'; -- increment address counter
				comp_value_int <= '1'; -- compare value
				reset_count_int <= '0';
         when others =>
            oe_n_int 	<= '1';
            we_n_int 	<= '1';
				dir_int 	<= '1'; -- read (output disabled)
				store_value_int <= '0';
				increment_int <= '0';
				comp_value_int <= '0';
				reset_count_int <= '1';
      end case;      
   end process;
 
   -- The Sram_test_next state Process is the combinatorial next
   -- state decode part of the Moore state machine 
   sram_test_next_state: process (state, count, start)
   begin
      next_state <= state;  --default is to stay in current state
      case (state) is
         when st1_w0_idle =>
			   -- run test one time on start condition
				if (start = '1') then
					next_state <= st2_w1_addr;
				else
					next_state <= st1_w0_idle;
				end if;
         when st2_w1_addr =>
            next_state <= st3_w2_data;
         when st3_w2_data =>
            next_state <= st4_w3_hold;
         when st4_w3_hold =>
            next_state <= st5_w4_d_en;
         when st5_w4_d_en =>
            next_state <= st6_w5_d_a;
         when st6_w5_d_a =>
			   -- goto read op if terminal count reached
            if (count = X"0003F") then --sim X"0003F", normal X"1FFFF"
					next_state <= st7_r0_idle;
				else
					next_state <= st2_w1_addr;
				end if;
         when st7_r0_idle =>
            next_state <= st8_r1_addr;
         when st8_r1_addr =>
            next_state <= st9_r2_oe;
         when st9_r2_oe =>
            next_state <= st10_r3_hold;
         when st10_r3_hold =>
            next_state <= st11_r4_data;
         when st11_r4_data =>
            next_state <= st12_r5_comp;
         when st12_r5_comp =>
			   -- test complete if terminal count reached
            if (count = X"0003F") then --sim X"0003F", normal X"1FFFF"
            	next_state <= st1_w0_idle; -- compare done
				else
					next_state <= st8_r1_addr;
				end if;
         when others =>
            next_state <= st1_w0_idle;
      end case;      
   end process;

   address_counter: process (sm_clk_in)
   begin
      if (sm_clk_in'event and sm_clk_in = '1') then
         if (rst_in = '1' or reset_count = '1') then
				count <= (others =>'0');
         else
				if (increment = '1') then
					count <= count + 1;
				else
					count <= count; --hold value
				end if;
         end if;        
      end if;
   end process;
	
   -- The Store Data process captures the data input value
	-- and the expected data (the address value) when instructed
	-- by the state machine.
   store_data: process (sm_clk_in)
   begin
      if (sm_clk_in'event and sm_clk_in = '1') then
         if (rst_in = '1') then
 				result <= (others =>'0');
				value <= (others =>'0');
         else
				if (store_value = '1') then
					value <= count(7 downto 0);
					result <= din;
				else
					value <= value; --hold value
					result <= result; --hold value
				end if;
         end if;        
      end if;
   end process;	
	
   -- The Error Counter process counts any errors that occur
   -- and creates an active high flag to indicate when any
   -- errors have been found. 	
   error_counter: process (sm_clk_in)
   begin
      if (sm_clk_in'event and sm_clk_in = '1') then
         if (start = '1') then
            errors_int 	<= (others =>'0');
				test_failed_int <= '0';
			else
				if (comp_value = '1') and (result /= value) then
					errors_int <= errors_int + 1;
					test_failed_int <= '1';
				else
					errors_int <= errors_int;
					test_failed_int <= test_failed_int;
				end if;
         end if;        
      end if;
   end process;

	-- connect internal signals to the port map
	errors <= errors_int;
	test_failed <= test_failed_int;
	a <= count;
	dout <= count(7 downto 0) when (dir_copy = '0') else X"00";

end rtl;

