`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:54:37 08/19/2013 
// Design Name: 
// Module Name:    Feistel_network 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Feistel_network(
    input [32:0] Input,
    output [32:0] Output,
    input encrypt_en
    );


endmodule
